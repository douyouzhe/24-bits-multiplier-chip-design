LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.all;
entity rom is
port(
ADDRESS: in std_logic_vector(16 downto 0);
ENA: in std_logic;
RD: in std_logic;
ROMINSTRUCTION:out std_logic_vector(23 downto 0)
);
end rom;
architecture ARCH of rom is
begin
process(ADDRESS,ENA,RD)
type rom_array is array(0 to 131055) of std_logic_vector(23 downto 0);
variable mem:rom_array:=( 
("000000000000000000000000"),
("000000000000000000000000"),
("000001000000000000000000"),
("000001100000000000000000"),
("111000000000000000000000"),
("000001100000000000000000"),
("111010000000000000000110"),
("111100000000000000000111"),
("101000000000000000001000"),
("000101000000000000000000"),
("110001100001010101010101"),
("000000000000000000000100"),
("111110000001010101010101"),
("110010000000000000000110"),
("000000000000000000000000"),
("000000000000000000000000"),
("000000000000000000000000"),
("000000000000000000000000"),
("000000000000000000000100"),
("000000000000000000000100"),
("000000000000000000000100"),
("000000000000000000000100"),
("000000000000000000000100"),
("000000000000000000000100"),
("000000000000000000000100"),
others=>("111111111111111111111111"));
begin
if(ENA='1' and RD='1')then
ROMINSTRUCTION<=mem((to_integer(unsigned(ADDRESS))));
else
ROMINSTRUCTION<=(others=>'Z');
end if;
end process;
end ARCH;